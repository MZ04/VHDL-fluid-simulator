----------------------------------------------------------------------------------
-- Team: LedMatrixGroup
-- Engineer: 
-- 
-- Create Date: 03/13/2025 04:43:41 PM
-- Module Name: display_driver - Behavioral
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity fsm is
--  Port ( );
end fsm;

architecture Behavioral of fsm is

begin


end Behavioral;
